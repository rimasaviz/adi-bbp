
module NCOTableLUT(
  input                                    clock,
  input      [9:0] addr,
  output reg [29:0] data
);
  always @(posedge clock) begin
    case (addr)
      10'b0: data <= 30'h0;
      10'b1: data <= 30'h1921fb;
      10'b10: data <= 30'h3243f1;
      10'b11: data <= 30'h4b65e1;
      10'b100: data <= 30'h6487c4;
      10'b101: data <= 30'h7da998;
      10'b110: data <= 30'h96cb58;
      10'b111: data <= 30'hafed02;
      10'b1000: data <= 30'hc90e90;
      10'b1001: data <= 30'he22fff;
      10'b1010: data <= 30'hfb514b;
      10'b1011: data <= 30'h1147271;
      10'b1100: data <= 30'h12d936c;
      10'b1101: data <= 30'h146b438;
      10'b1110: data <= 30'h15fd4d2;
      10'b1111: data <= 30'h178f536;
      10'b10000: data <= 30'h192155f;
      10'b10001: data <= 30'h1ab354b;
      10'b10010: data <= 30'h1c454f5;
      10'b10011: data <= 30'h1dd7459;
      10'b10100: data <= 30'h1f69373;
      10'b10101: data <= 30'h20fb240;
      10'b10110: data <= 30'h228d0bb;
      10'b10111: data <= 30'h241eee2;
      10'b11000: data <= 30'h25b0caf;
      10'b11001: data <= 30'h2742a1f;
      10'b11010: data <= 30'h28d472e;
      10'b11011: data <= 30'h2a663d8;
      10'b11100: data <= 30'h2bf801a;
      10'b11101: data <= 30'h2d89bf0;
      10'b11110: data <= 30'h2f1b755;
      10'b11111: data <= 30'h30ad245;
      10'b100000: data <= 30'h323ecbe;
      10'b100001: data <= 30'h33d06bb;
      10'b100010: data <= 30'h3562038;
      10'b100011: data <= 30'h36f3931;
      10'b100100: data <= 30'h38851a2;
      10'b100101: data <= 30'h3a16988;
      10'b100110: data <= 30'h3ba80df;
      10'b100111: data <= 30'h3d397a3;
      10'b101000: data <= 30'h3ecadcf;
      10'b101001: data <= 30'h405c361;
      10'b101010: data <= 30'h41ed854;
      10'b101011: data <= 30'h437eca4;
      10'b101100: data <= 30'h451004d;
      10'b101101: data <= 30'h46a134c;
      10'b101110: data <= 30'h483259d;
      10'b101111: data <= 30'h49c373c;
      10'b110000: data <= 30'h4b54825;
      10'b110001: data <= 30'h4ce5854;
      10'b110010: data <= 30'h4e767c5;
      10'b110011: data <= 30'h5007674;
      10'b110100: data <= 30'h519845e;
      10'b110101: data <= 30'h532917f;
      10'b110110: data <= 30'h54b9dd3;
      10'b110111: data <= 30'h564a955;
      10'b111000: data <= 30'h57db403;
      10'b111001: data <= 30'h596bdd7;
      10'b111010: data <= 30'h5afc6d0;
      10'b111011: data <= 30'h5c8cee7;
      10'b111100: data <= 30'h5e1d61b;
      10'b111101: data <= 30'h5fadc66;
      10'b111110: data <= 30'h613e1c5;
      10'b111111: data <= 30'h62ce634;
      10'b1000000: data <= 30'h645e9af;
      10'b1000001: data <= 30'h65eec33;
      10'b1000010: data <= 30'h677edbb;
      10'b1000011: data <= 30'h690ee44;
      10'b1000100: data <= 30'h6a9edc9;
      10'b1000101: data <= 30'h6c2ec48;
      10'b1000110: data <= 30'h6dbe9bb;
      10'b1000111: data <= 30'h6f4e620;
      10'b1001000: data <= 30'h70de172;
      10'b1001001: data <= 30'h726dbae;
      10'b1001010: data <= 30'h73fd4cf;
      10'b1001011: data <= 30'h758ccd2;
      10'b1001100: data <= 30'h771c3b3;
      10'b1001101: data <= 30'h78ab96e;
      10'b1001110: data <= 30'h7a3adff;
      10'b1001111: data <= 30'h7bca163;
      10'b1010000: data <= 30'h7d59396;
      10'b1010001: data <= 30'h7ee8493;
      10'b1010010: data <= 30'h8077457;
      10'b1010011: data <= 30'h82062de;
      10'b1010100: data <= 30'h8395024;
      10'b1010101: data <= 30'h8523c25;
      10'b1010110: data <= 30'h86b26de;
      10'b1010111: data <= 30'h884104b;
      10'b1011000: data <= 30'h89cf867;
      10'b1011001: data <= 30'h8b5df30;
      10'b1011010: data <= 30'h8cec4a0;
      10'b1011011: data <= 30'h8e7a8b5;
      10'b1011100: data <= 30'h9008b6a;
      10'b1011101: data <= 30'h9196cbc;
      10'b1011110: data <= 30'h9324ca7;
      10'b1011111: data <= 30'h94b2b27;
      10'b1100000: data <= 30'h9640837;
      10'b1100001: data <= 30'h97ce3d5;
      10'b1100010: data <= 30'h995bdfd;
      10'b1100011: data <= 30'h9ae96aa;
      10'b1100100: data <= 30'h9c76dd8;
      10'b1100101: data <= 30'h9e04385;
      10'b1100110: data <= 30'h9f917ac;
      10'b1100111: data <= 30'ha11ea49;
      10'b1101000: data <= 30'ha2abb59;
      10'b1101001: data <= 30'ha438ad7;
      10'b1101010: data <= 30'ha5c58c0;
      10'b1101011: data <= 30'ha752510;
      10'b1101100: data <= 30'ha8defc3;
      10'b1101101: data <= 30'haa6b8d5;
      10'b1101110: data <= 30'habf8043;
      10'b1101111: data <= 30'had84609;
      10'b1110000: data <= 30'haf10a22;
      10'b1110001: data <= 30'hb09cc8c;
      10'b1110010: data <= 30'hb228d42;
      10'b1110011: data <= 30'hb3b4c40;
      10'b1110100: data <= 30'hb540982;
      10'b1110101: data <= 30'hb6cc506;
      10'b1110110: data <= 30'hb857ec7;
      10'b1110111: data <= 30'hb9e36c0;
      10'b1111000: data <= 30'hbb6ecef;
      10'b1111001: data <= 30'hbcfa150;
      10'b1111010: data <= 30'hbe853de;
      10'b1111011: data <= 30'hc010496;
      10'b1111100: data <= 30'hc19b374;
      10'b1111101: data <= 30'hc326075;
      10'b1111110: data <= 30'hc4b0b94;
      10'b1111111: data <= 30'hc63b4ce;
      10'b10000000: data <= 30'hc7c5c1e;
      10'b10000001: data <= 30'hc950182;
      10'b10000010: data <= 30'hcada4f5;
      10'b10000011: data <= 30'hcc64673;
      10'b10000100: data <= 30'hcdee5f9;
      10'b10000101: data <= 30'hcf78383;
      10'b10000110: data <= 30'hd101f0e;
      10'b10000111: data <= 30'hd28b894;
      10'b10001000: data <= 30'hd415013;
      10'b10001001: data <= 30'hd59e586;
      10'b10001010: data <= 30'hd7278eb;
      10'b10001011: data <= 30'hd8b0a3d;
      10'b10001100: data <= 30'hda39978;
      10'b10001101: data <= 30'hdbc2698;
      10'b10001110: data <= 30'hdd4b19a;
      10'b10001111: data <= 30'hded3a7b;
      10'b10010000: data <= 30'he05c135;
      10'b10010001: data <= 30'he1e45c6;
      10'b10010010: data <= 30'he36c82a;
      10'b10010011: data <= 30'he4f485c;
      10'b10010100: data <= 30'he67c65a;
      10'b10010101: data <= 30'he80421e;
      10'b10010110: data <= 30'he98bba7;
      10'b10010111: data <= 30'heb132ef;
      10'b10011000: data <= 30'hec9a7f3;
      10'b10011001: data <= 30'hee21aaf;
      10'b10011010: data <= 30'hefa8b20;
      10'b10011011: data <= 30'hf12f941;
      10'b10011100: data <= 30'hf2b650f;
      10'b10011101: data <= 30'hf43ce86;
      10'b10011110: data <= 30'hf5c35a3;
      10'b10011111: data <= 30'hf749a61;
      10'b10100000: data <= 30'hf8cfcbe;
      10'b10100001: data <= 30'hfa55cb4;
      10'b10100010: data <= 30'hfbdba40;
      10'b10100011: data <= 30'hfd6155f;
      10'b10100100: data <= 30'hfee6e0d;
      10'b10100101: data <= 30'h1006c446;
      10'b10100110: data <= 30'h101f1807;
      10'b10100111: data <= 30'h1037694b;
      10'b10101000: data <= 30'h104fb80e;
      10'b10101001: data <= 30'h1068044e;
      10'b10101010: data <= 30'h10804e06;
      10'b10101011: data <= 30'h10989532;
      10'b10101100: data <= 30'h10b0d9d0;
      10'b10101101: data <= 30'h10c91bda;
      10'b10101110: data <= 30'h10e15b4e;
      10'b10101111: data <= 30'h10f99827;
      10'b10110000: data <= 30'h1111d263;
      10'b10110001: data <= 30'h112a09fc;
      10'b10110010: data <= 30'h11423ef0;
      10'b10110011: data <= 30'h115a713a;
      10'b10110100: data <= 30'h1172a0d7;
      10'b10110101: data <= 30'h118acdc4;
      10'b10110110: data <= 30'h11a2f7fc;
      10'b10110111: data <= 30'h11bb1f7c;
      10'b10111000: data <= 30'h11d3443f;
      10'b10111001: data <= 30'h11eb6643;
      10'b10111010: data <= 30'h12038584;
      10'b10111011: data <= 30'h121ba1fd;
      10'b10111100: data <= 30'h1233bbac;
      10'b10111101: data <= 30'h124bd28c;
      10'b10111110: data <= 30'h1263e699;
      10'b10111111: data <= 30'h127bf7d1;
      10'b11000000: data <= 30'h1294062f;
      10'b11000001: data <= 30'h12ac11af;
      10'b11000010: data <= 30'h12c41a4f;
      10'b11000011: data <= 30'h12dc2009;
      10'b11000100: data <= 30'h12f422db;
      10'b11000101: data <= 30'h130c22c1;
      10'b11000110: data <= 30'h13241fb6;
      10'b11000111: data <= 30'h133c19b8;
      10'b11001000: data <= 30'h135410c3;
      10'b11001001: data <= 30'h136c04d2;
      10'b11001010: data <= 30'h1383f5e3;
      10'b11001011: data <= 30'h139be3f2;
      10'b11001100: data <= 30'h13b3cefa;
      10'b11001101: data <= 30'h13cbb6f8;
      10'b11001110: data <= 30'h13e39be9;
      10'b11001111: data <= 30'h13fb7dc9;
      10'b11010000: data <= 30'h14135c94;
      10'b11010001: data <= 30'h142b3846;
      10'b11010010: data <= 30'h144310dd;
      10'b11010011: data <= 30'h145ae653;
      10'b11010100: data <= 30'h1472b8a5;
      10'b11010101: data <= 30'h148a87d1;
      10'b11010110: data <= 30'h14a253d1;
      10'b11010111: data <= 30'h14ba1ca3;
      10'b11011000: data <= 30'h14d1e242;
      10'b11011001: data <= 30'h14e9a4ac;
      10'b11011010: data <= 30'h150163dc;
      10'b11011011: data <= 30'h15191fcf;
      10'b11011100: data <= 30'h1530d881;
      10'b11011101: data <= 30'h15488dee;
      10'b11011110: data <= 30'h15604013;
      10'b11011111: data <= 30'h1577eeec;
      10'b11100000: data <= 30'h158f9a76;
      10'b11100001: data <= 30'h15a742ac;
      10'b11100010: data <= 30'h15bee78c;
      10'b11100011: data <= 30'h15d68911;
      10'b11100100: data <= 30'h15ee2738;
      10'b11100101: data <= 30'h1605c1fd;
      10'b11100110: data <= 30'h161d595d;
      10'b11100111: data <= 30'h1634ed53;
      10'b11101000: data <= 30'h164c7ddd;
      10'b11101001: data <= 30'h16640af7;
      10'b11101010: data <= 30'h167b949d;
      10'b11101011: data <= 30'h16931acb;
      10'b11101100: data <= 30'h16aa9d7e;
      10'b11101101: data <= 30'h16c21cb2;
      10'b11101110: data <= 30'h16d99864;
      10'b11101111: data <= 30'h16f1108f;
      10'b11110000: data <= 30'h17088531;
      10'b11110001: data <= 30'h171ff646;
      10'b11110010: data <= 30'h173763c9;
      10'b11110011: data <= 30'h174ecdb8;
      10'b11110100: data <= 30'h1766340f;
      10'b11110101: data <= 30'h177d96ca;
      10'b11110110: data <= 30'h1794f5e6;
      10'b11110111: data <= 30'h17ac515f;
      10'b11111000: data <= 30'h17c3a931;
      10'b11111001: data <= 30'h17dafd59;
      10'b11111010: data <= 30'h17f24dd3;
      10'b11111011: data <= 30'h18099a9c;
      10'b11111100: data <= 30'h1820e3b0;
      10'b11111101: data <= 30'h1838290c;
      10'b11111110: data <= 30'h184f6aab;
      10'b11111111: data <= 30'h1866a88a;
      10'b100000000: data <= 30'h187de2a7;
      10'b100000001: data <= 30'h189518fc;
      10'b100000010: data <= 30'h18ac4b87;
      10'b100000011: data <= 30'h18c37a44;
      10'b100000100: data <= 30'h18daa52f;
      10'b100000101: data <= 30'h18f1cc45;
      10'b100000110: data <= 30'h1908ef82;
      10'b100000111: data <= 30'h19200ee3;
      10'b100001000: data <= 30'h19372a64;
      10'b100001001: data <= 30'h194e4201;
      10'b100001010: data <= 30'h196555b8;
      10'b100001011: data <= 30'h197c6584;
      10'b100001100: data <= 30'h19937161;
      10'b100001101: data <= 30'h19aa794d;
      10'b100001110: data <= 30'h19c17d44;
      10'b100001111: data <= 30'h19d87d42;
      10'b100010000: data <= 30'h19ef7944;
      10'b100010001: data <= 30'h1a067145;
      10'b100010010: data <= 30'h1a1d6544;
      10'b100010011: data <= 30'h1a34553b;
      10'b100010100: data <= 30'h1a4b4128;
      10'b100010101: data <= 30'h1a622907;
      10'b100010110: data <= 30'h1a790cd4;
      10'b100010111: data <= 30'h1a8fec8c;
      10'b100011000: data <= 30'h1aa6c82b;
      10'b100011001: data <= 30'h1abd9faf;
      10'b100011010: data <= 30'h1ad47312;
      10'b100011011: data <= 30'h1aeb4253;
      10'b100011100: data <= 30'h1b020d6c;
      10'b100011101: data <= 30'h1b18d45c;
      10'b100011110: data <= 30'h1b2f971e;
      10'b100011111: data <= 30'h1b4655ae;
      10'b100100000: data <= 30'h1b5d100a;
      10'b100100001: data <= 30'h1b73c62d;
      10'b100100010: data <= 30'h1b8a7815;
      10'b100100011: data <= 30'h1ba125bd;
      10'b100100100: data <= 30'h1bb7cf23;
      10'b100100101: data <= 30'h1bce7442;
      10'b100100110: data <= 30'h1be51518;
      10'b100100111: data <= 30'h1bfbb1a0;
      10'b100101000: data <= 30'h1c1249d8;
      10'b100101001: data <= 30'h1c28ddbb;
      10'b100101010: data <= 30'h1c3f6d47;
      10'b100101011: data <= 30'h1c55f878;
      10'b100101100: data <= 30'h1c6c7f4a;
      10'b100101101: data <= 30'h1c8301b9;
      10'b100101110: data <= 30'h1c997fc4;
      10'b100101111: data <= 30'h1caff965;
      10'b100110000: data <= 30'h1cc66e99;
      10'b100110001: data <= 30'h1cdcdf5e;
      10'b100110010: data <= 30'h1cf34baf;
      10'b100110011: data <= 30'h1d09b389;
      10'b100110100: data <= 30'h1d2016e9;
      10'b100110101: data <= 30'h1d3675cb;
      10'b100110110: data <= 30'h1d4cd02c;
      10'b100110111: data <= 30'h1d632608;
      10'b100111000: data <= 30'h1d79775c;
      10'b100111001: data <= 30'h1d8fc424;
      10'b100111010: data <= 30'h1da60c5d;
      10'b100111011: data <= 30'h1dbc5004;
      10'b100111100: data <= 30'h1dd28f15;
      10'b100111101: data <= 30'h1de8c98c;
      10'b100111110: data <= 30'h1dfeff67;
      10'b100111111: data <= 30'h1e1530a1;
      10'b101000000: data <= 30'h1e2b5d38;
      10'b101000001: data <= 30'h1e418528;
      10'b101000010: data <= 30'h1e57a86d;
      10'b101000011: data <= 30'h1e6dc705;
      10'b101000100: data <= 30'h1e83e0eb;
      10'b101000101: data <= 30'h1e99f61d;
      10'b101000110: data <= 30'h1eb00696;
      10'b101000111: data <= 30'h1ec61254;
      10'b101001000: data <= 30'h1edc1953;
      10'b101001001: data <= 30'h1ef21b90;
      10'b101001010: data <= 30'h1f081907;
      10'b101001011: data <= 30'h1f1e11b5;
      10'b101001100: data <= 30'h1f340596;
      10'b101001101: data <= 30'h1f49f4a8;
      10'b101001110: data <= 30'h1f5fdee6;
      10'b101001111: data <= 30'h1f75c44e;
      10'b101010000: data <= 30'h1f8ba4dc;
      10'b101010001: data <= 30'h1fa1808c;
      10'b101010010: data <= 30'h1fb7575c;
      10'b101010011: data <= 30'h1fcd2948;
      10'b101010100: data <= 30'h1fe2f64c;
      10'b101010101: data <= 30'h1ff8be65;
      10'b101010110: data <= 30'h200e8190;
      10'b101010111: data <= 30'h20243fca;
      10'b101011000: data <= 30'h2039f90f;
      10'b101011001: data <= 30'h204fad5b;
      10'b101011010: data <= 30'h20655cac;
      10'b101011011: data <= 30'h207b06fe;
      10'b101011100: data <= 30'h2090ac4d;
      10'b101011101: data <= 30'h20a64c97;
      10'b101011110: data <= 30'h20bbe7d8;
      10'b101011111: data <= 30'h20d17e0d;
      10'b101100000: data <= 30'h20e70f32;
      10'b101100001: data <= 30'h20fc9b44;
      10'b101100010: data <= 30'h21122240;
      10'b101100011: data <= 30'h2127a423;
      10'b101100100: data <= 30'h213d20e8;
      10'b101100101: data <= 30'h2152988d;
      10'b101100110: data <= 30'h21680b0f;
      10'b101100111: data <= 30'h217d786a;
      10'b101101000: data <= 30'h2192e09b;
      10'b101101001: data <= 30'h21a8439e;
      10'b101101010: data <= 30'h21bda171;
      10'b101101011: data <= 30'h21d2fa0f;
      10'b101101100: data <= 30'h21e84d76;
      10'b101101101: data <= 30'h21fd9ba3;
      10'b101101110: data <= 30'h2212e492;
      10'b101101111: data <= 30'h2228283f;
      10'b101110000: data <= 30'h223d66a8;
      10'b101110001: data <= 30'h22529fca;
      10'b101110010: data <= 30'h2267d3a0;
      10'b101110011: data <= 30'h227d0228;
      10'b101110100: data <= 30'h22922b5e;
      10'b101110101: data <= 30'h22a74f40;
      10'b101110110: data <= 30'h22bc6dca;
      10'b101110111: data <= 30'h22d186f8;
      10'b101111000: data <= 30'h22e69ac8;
      10'b101111001: data <= 30'h22fba936;
      10'b101111010: data <= 30'h2310b23e;
      10'b101111011: data <= 30'h2325b5df;
      10'b101111100: data <= 30'h233ab414;
      10'b101111101: data <= 30'h234facda;
      10'b101111110: data <= 30'h2364a02e;
      10'b101111111: data <= 30'h23798e0d;
      10'b110000000: data <= 30'h238e7673;
      10'b110000001: data <= 30'h23a3595e;
      10'b110000010: data <= 30'h23b836ca;
      10'b110000011: data <= 30'h23cd0eb3;
      10'b110000100: data <= 30'h23e1e117;
      10'b110000101: data <= 30'h23f6adf3;
      10'b110000110: data <= 30'h240b7543;
      10'b110000111: data <= 30'h24203704;
      10'b110001000: data <= 30'h2434f332;
      10'b110001001: data <= 30'h2449a9cc;
      10'b110001010: data <= 30'h245e5acc;
      10'b110001011: data <= 30'h24730631;
      10'b110001100: data <= 30'h2487abf7;
      10'b110001101: data <= 30'h249c4c1b;
      10'b110001110: data <= 30'h24b0e699;
      10'b110001111: data <= 30'h24c57b6f;
      10'b110010000: data <= 30'h24da0a9a;
      10'b110010001: data <= 30'h24ee9415;
      10'b110010010: data <= 30'h250317df;
      10'b110010011: data <= 30'h251795f3;
      10'b110010100: data <= 30'h252c0e4f;
      10'b110010101: data <= 30'h254080ef;
      10'b110010110: data <= 30'h2554edd1;
      10'b110010111: data <= 30'h256954f1;
      10'b110011000: data <= 30'h257db64c;
      10'b110011001: data <= 30'h259211df;
      10'b110011010: data <= 30'h25a667a7;
      10'b110011011: data <= 30'h25bab7a0;
      10'b110011100: data <= 30'h25cf01c8;
      10'b110011101: data <= 30'h25e3461b;
      10'b110011110: data <= 30'h25f78497;
      10'b110011111: data <= 30'h260bbd37;
      10'b110100000: data <= 30'h261feffa;
      10'b110100001: data <= 30'h26341cdb;
      10'b110100010: data <= 30'h264843d9;
      10'b110100011: data <= 30'h265c64ef;
      10'b110100100: data <= 30'h2670801a;
      10'b110100101: data <= 30'h26849558;
      10'b110100110: data <= 30'h2698a4a6;
      10'b110100111: data <= 30'h26acadff;
      10'b110101000: data <= 30'h26c0b162;
      10'b110101001: data <= 30'h26d4aecb;
      10'b110101010: data <= 30'h26e8a637;
      10'b110101011: data <= 30'h26fc97a3;
      10'b110101100: data <= 30'h2710830c;
      10'b110101101: data <= 30'h2724686e;
      10'b110101110: data <= 30'h273847c8;
      10'b110101111: data <= 30'h274c2115;
      10'b110110000: data <= 30'h275ff452;
      10'b110110001: data <= 30'h2773c17d;
      10'b110110010: data <= 30'h27878893;
      10'b110110011: data <= 30'h279b4990;
      10'b110110100: data <= 30'h27af0472;
      10'b110110101: data <= 30'h27c2b934;
      10'b110110110: data <= 30'h27d667d5;
      10'b110110111: data <= 30'h27ea1052;
      10'b110111000: data <= 30'h27fdb2a7;
      10'b110111001: data <= 30'h28114ed0;
      10'b110111010: data <= 30'h2824e4cc;
      10'b110111011: data <= 30'h28387498;
      10'b110111100: data <= 30'h284bfe2f;
      10'b110111101: data <= 30'h285f8190;
      10'b110111110: data <= 30'h2872feb6;
      10'b110111111: data <= 30'h288675a0;
      10'b111000000: data <= 30'h2899e64a;
      10'b111000001: data <= 30'h28ad50b1;
      10'b111000010: data <= 30'h28c0b4d2;
      10'b111000011: data <= 30'h28d412ab;
      10'b111000100: data <= 30'h28e76a37;
      10'b111000101: data <= 30'h28fabb75;
      10'b111000110: data <= 30'h290e0661;
      10'b111000111: data <= 30'h29214af8;
      10'b111001000: data <= 30'h29348937;
      10'b111001001: data <= 30'h2947c11c;
      10'b111001010: data <= 30'h295af2a3;
      10'b111001011: data <= 30'h296e1dc9;
      10'b111001100: data <= 30'h2981428c;
      10'b111001101: data <= 30'h299460e8;
      10'b111001110: data <= 30'h29a778db;
      10'b111001111: data <= 30'h29ba8a61;
      10'b111010000: data <= 30'h29cd9578;
      10'b111010001: data <= 30'h29e09a1c;
      10'b111010010: data <= 30'h29f3984c;
      10'b111010011: data <= 30'h2a069003;
      10'b111010100: data <= 30'h2a19813f;
      10'b111010101: data <= 30'h2a2c6bfd;
      10'b111010110: data <= 30'h2a3f503a;
      10'b111010111: data <= 30'h2a522df3;
      10'b111011000: data <= 30'h2a650525;
      10'b111011001: data <= 30'h2a77d5ce;
      10'b111011010: data <= 30'h2a8a9fea;
      10'b111011011: data <= 30'h2a9d6377;
      10'b111011100: data <= 30'h2ab02071;
      10'b111011101: data <= 30'h2ac2d6d6;
      10'b111011110: data <= 30'h2ad586a3;
      10'b111011111: data <= 30'h2ae82fd5;
      10'b111100000: data <= 30'h2afad269;
      10'b111100001: data <= 30'h2b0d6e5c;
      10'b111100010: data <= 30'h2b2003ac;
      10'b111100011: data <= 30'h2b329255;
      10'b111100100: data <= 30'h2b451a55;
      10'b111100101: data <= 30'h2b579ba8;
      10'b111100110: data <= 30'h2b6a164d;
      10'b111100111: data <= 30'h2b7c8a3f;
      10'b111101000: data <= 30'h2b8ef77d;
      10'b111101001: data <= 30'h2ba15e03;
      10'b111101010: data <= 30'h2bb3bdce;
      10'b111101011: data <= 30'h2bc616dd;
      10'b111101100: data <= 30'h2bd8692b;
      10'b111101101: data <= 30'h2beab4b6;
      10'b111101110: data <= 30'h2bfcf97c;
      10'b111101111: data <= 30'h2c0f3779;
      10'b111110000: data <= 30'h2c216eaa;
      10'b111110001: data <= 30'h2c339f0e;
      10'b111110010: data <= 30'h2c45c8a0;
      10'b111110011: data <= 30'h2c57eb5e;
      10'b111110100: data <= 30'h2c6a0746;
      10'b111110101: data <= 30'h2c7c1c55;
      10'b111110110: data <= 30'h2c8e2a87;
      10'b111110111: data <= 30'h2ca031da;
      10'b111111000: data <= 30'h2cb2324c;
      10'b111111001: data <= 30'h2cc42bd9;
      10'b111111010: data <= 30'h2cd61e7f;
      10'b111111011: data <= 30'h2ce80a3a;
      10'b111111100: data <= 30'h2cf9ef09;
      10'b111111101: data <= 30'h2d0bcce8;
      10'b111111110: data <= 30'h2d1da3d5;
      10'b111111111: data <= 30'h2d2f73cd;
      10'b1000000000: data <= 30'h2d413ccd;
      10'b1000000001: data <= 30'h2d52fed2;
      10'b1000000010: data <= 30'h2d64b9da;
      10'b1000000011: data <= 30'h2d766de2;
      10'b1000000100: data <= 30'h2d881ae8;
      10'b1000000101: data <= 30'h2d99c0e7;
      10'b1000000110: data <= 30'h2dab5fdf;
      10'b1000000111: data <= 30'h2dbcf7cb;
      10'b1000001000: data <= 30'h2dce88aa;
      10'b1000001001: data <= 30'h2de01278;
      10'b1000001010: data <= 30'h2df19534;
      10'b1000001011: data <= 30'h2e0310d9;
      10'b1000001100: data <= 30'h2e148566;
      10'b1000001101: data <= 30'h2e25f2d8;
      10'b1000001110: data <= 30'h2e37592c;
      10'b1000001111: data <= 30'h2e48b860;
      10'b1000010000: data <= 30'h2e5a1070;
      10'b1000010001: data <= 30'h2e6b615a;
      10'b1000010010: data <= 30'h2e7cab1c;
      10'b1000010011: data <= 30'h2e8dedb3;
      10'b1000010100: data <= 30'h2e9f291b;
      10'b1000010101: data <= 30'h2eb05d53;
      10'b1000010110: data <= 30'h2ec18a58;
      10'b1000010111: data <= 30'h2ed2b027;
      10'b1000011000: data <= 30'h2ee3cebe;
      10'b1000011001: data <= 30'h2ef4e619;
      10'b1000011010: data <= 30'h2f05f637;
      10'b1000011011: data <= 30'h2f16ff14;
      10'b1000011100: data <= 30'h2f2800af;
      10'b1000011101: data <= 30'h2f38fb03;
      10'b1000011110: data <= 30'h2f49ee0f;
      10'b1000011111: data <= 30'h2f5ad9d1;
      10'b1000100000: data <= 30'h2f6bbe45;
      10'b1000100001: data <= 30'h2f7c9b69;
      10'b1000100010: data <= 30'h2f8d713a;
      10'b1000100011: data <= 30'h2f9e3fb6;
      10'b1000100100: data <= 30'h2faf06da;
      10'b1000100101: data <= 30'h2fbfc6a3;
      10'b1000100110: data <= 30'h2fd07f0f;
      10'b1000100111: data <= 30'h2fe1301c;
      10'b1000101000: data <= 30'h2ff1d9c7;
      10'b1000101001: data <= 30'h30027c0c;
      10'b1000101010: data <= 30'h301316eb;
      10'b1000101011: data <= 30'h3023aa5f;
      10'b1000101100: data <= 30'h30343667;
      10'b1000101101: data <= 30'h3044bb00;
      10'b1000101110: data <= 30'h30553828;
      10'b1000101111: data <= 30'h3065addb;
      10'b1000110000: data <= 30'h30761c18;
      10'b1000110001: data <= 30'h308682dc;
      10'b1000110010: data <= 30'h3096e223;
      10'b1000110011: data <= 30'h30a739ed;
      10'b1000110100: data <= 30'h30b78a36;
      10'b1000110101: data <= 30'h30c7d2fb;
      10'b1000110110: data <= 30'h30d8143b;
      10'b1000110111: data <= 30'h30e84df3;
      10'b1000111000: data <= 30'h30f8801f;
      10'b1000111001: data <= 30'h3108aabf;
      10'b1000111010: data <= 30'h3118cdcf;
      10'b1000111011: data <= 30'h3128e94c;
      10'b1000111100: data <= 30'h3138fd35;
      10'b1000111101: data <= 30'h31490986;
      10'b1000111110: data <= 30'h31590e3e;
      10'b1000111111: data <= 30'h31690b59;
      10'b1001000000: data <= 30'h317900d6;
      10'b1001000001: data <= 30'h3188eeb2;
      10'b1001000010: data <= 30'h3198d4ea;
      10'b1001000011: data <= 30'h31a8b37c;
      10'b1001000100: data <= 30'h31b88a66;
      10'b1001000101: data <= 30'h31c859a5;
      10'b1001000110: data <= 30'h31d82137;
      10'b1001000111: data <= 30'h31e7e118;
      10'b1001001000: data <= 30'h31f79948;
      10'b1001001001: data <= 30'h320749c3;
      10'b1001001010: data <= 30'h3216f287;
      10'b1001001011: data <= 30'h32269391;
      10'b1001001100: data <= 30'h32362ce0;
      10'b1001001101: data <= 30'h3245be70;
      10'b1001001110: data <= 30'h32554840;
      10'b1001001111: data <= 30'h3264ca4c;
      10'b1001010000: data <= 30'h32744493;
      10'b1001010001: data <= 30'h3283b712;
      10'b1001010010: data <= 30'h329321c7;
      10'b1001010011: data <= 30'h32a284b0;
      10'b1001010100: data <= 30'h32b1dfc9;
      10'b1001010101: data <= 30'h32c13311;
      10'b1001010110: data <= 30'h32d07e85;
      10'b1001010111: data <= 30'h32dfc224;
      10'b1001011000: data <= 30'h32eefdea;
      10'b1001011001: data <= 30'h32fe31d5;
      10'b1001011010: data <= 30'h330d5de3;
      10'b1001011011: data <= 30'h331c8211;
      10'b1001011100: data <= 30'h332b9e5e;
      10'b1001011101: data <= 30'h333ab2c6;
      10'b1001011110: data <= 30'h3349bf48;
      10'b1001011111: data <= 30'h3358c3e2;
      10'b1001100000: data <= 30'h3367c090;
      10'b1001100001: data <= 30'h3376b551;
      10'b1001100010: data <= 30'h3385a222;
      10'b1001100011: data <= 30'h33948701;
      10'b1001100100: data <= 30'h33a363ec;
      10'b1001100101: data <= 30'h33b238e0;
      10'b1001100110: data <= 30'h33c105db;
      10'b1001100111: data <= 30'h33cfcadc;
      10'b1001101000: data <= 30'h33de87de;
      10'b1001101001: data <= 30'h33ed3ce1;
      10'b1001101010: data <= 30'h33fbe9e2;
      10'b1001101011: data <= 30'h340a8edf;
      10'b1001101100: data <= 30'h34192bd5;
      10'b1001101101: data <= 30'h3427c0c3;
      10'b1001101110: data <= 30'h34364da6;
      10'b1001101111: data <= 30'h3444d27b;
      10'b1001110000: data <= 30'h34534f41;
      10'b1001110001: data <= 30'h3461c3f5;
      10'b1001110010: data <= 30'h34703095;
      10'b1001110011: data <= 30'h347e951f;
      10'b1001110100: data <= 30'h348cf190;
      10'b1001110101: data <= 30'h349b45e7;
      10'b1001110110: data <= 30'h34a99221;
      10'b1001110111: data <= 30'h34b7d63c;
      10'b1001111000: data <= 30'h34c61236;
      10'b1001111001: data <= 30'h34d4460c;
      10'b1001111010: data <= 30'h34e271bd;
      10'b1001111011: data <= 30'h34f09546;
      10'b1001111100: data <= 30'h34feb0a5;
      10'b1001111101: data <= 30'h350cc3d8;
      10'b1001111110: data <= 30'h351acedd;
      10'b1001111111: data <= 30'h3528d1b1;
      10'b1010000000: data <= 30'h3536cc52;
      10'b1010000001: data <= 30'h3544bebf;
      10'b1010000010: data <= 30'h3552a8f4;
      10'b1010000011: data <= 30'h35608af1;
      10'b1010000100: data <= 30'h356e64b2;
      10'b1010000101: data <= 30'h357c3636;
      10'b1010000110: data <= 30'h3589ff7a;
      10'b1010000111: data <= 30'h3597c07d;
      10'b1010001000: data <= 30'h35a5793c;
      10'b1010001001: data <= 30'h35b329b5;
      10'b1010001010: data <= 30'h35c0d1e7;
      10'b1010001011: data <= 30'h35ce71ce;
      10'b1010001100: data <= 30'h35dc0968;
      10'b1010001101: data <= 30'h35e998b5;
      10'b1010001110: data <= 30'h35f71fb1;
      10'b1010001111: data <= 30'h36049e5b;
      10'b1010010000: data <= 30'h361214b0;
      10'b1010010001: data <= 30'h361f82af;
      10'b1010010010: data <= 30'h362ce855;
      10'b1010010011: data <= 30'h363a45a0;
      10'b1010010100: data <= 30'h36479a8e;
      10'b1010010101: data <= 30'h3654e71d;
      10'b1010010110: data <= 30'h36622b4c;
      10'b1010010111: data <= 30'h366f6717;
      10'b1010011000: data <= 30'h367c9a7e;
      10'b1010011001: data <= 30'h3689c57d;
      10'b1010011010: data <= 30'h3696e814;
      10'b1010011011: data <= 30'h36a4023f;
      10'b1010011100: data <= 30'h36b113fd;
      10'b1010011101: data <= 30'h36be1d4c;
      10'b1010011110: data <= 30'h36cb1e2a;
      10'b1010011111: data <= 30'h36d81695;
      10'b1010100000: data <= 30'h36e5068a;
      10'b1010100001: data <= 30'h36f1ee09;
      10'b1010100010: data <= 30'h36fecd0e;
      10'b1010100011: data <= 30'h370ba398;
      10'b1010100100: data <= 30'h371871a5;
      10'b1010100101: data <= 30'h37253733;
      10'b1010100110: data <= 30'h3731f440;
      10'b1010100111: data <= 30'h373ea8ca;
      10'b1010101000: data <= 30'h374b54ce;
      10'b1010101001: data <= 30'h3757f84c;
      10'b1010101010: data <= 30'h37649341;
      10'b1010101011: data <= 30'h377125ac;
      10'b1010101100: data <= 30'h377daf89;
      10'b1010101101: data <= 30'h378a30d8;
      10'b1010101110: data <= 30'h3796a996;
      10'b1010101111: data <= 30'h37a319c2;
      10'b1010110000: data <= 30'h37af8159;
      10'b1010110001: data <= 30'h37bbe05a;
      10'b1010110010: data <= 30'h37c836c2;
      10'b1010110011: data <= 30'h37d48490;
      10'b1010110100: data <= 30'h37e0c9c3;
      10'b1010110101: data <= 30'h37ed0657;
      10'b1010110110: data <= 30'h37f93a4b;
      10'b1010110111: data <= 30'h3805659e;
      10'b1010111000: data <= 30'h3811884d;
      10'b1010111001: data <= 30'h381da256;
      10'b1010111010: data <= 30'h3829b3b9;
      10'b1010111011: data <= 30'h3835bc71;
      10'b1010111100: data <= 30'h3841bc7f;
      10'b1010111101: data <= 30'h384db3e0;
      10'b1010111110: data <= 30'h3859a292;
      10'b1010111111: data <= 30'h38658894;
      10'b1011000000: data <= 30'h387165e3;
      10'b1011000001: data <= 30'h387d3a7e;
      10'b1011000010: data <= 30'h38890663;
      10'b1011000011: data <= 30'h3894c98f;
      10'b1011000100: data <= 30'h38a08402;
      10'b1011000101: data <= 30'h38ac35ba;
      10'b1011000110: data <= 30'h38b7deb4;
      10'b1011000111: data <= 30'h38c37eef;
      10'b1011001000: data <= 30'h38cf1669;
      10'b1011001001: data <= 30'h38daa520;
      10'b1011001010: data <= 30'h38e62b13;
      10'b1011001011: data <= 30'h38f1a840;
      10'b1011001100: data <= 30'h38fd1ca4;
      10'b1011001101: data <= 30'h3908883f;
      10'b1011001110: data <= 30'h3913eb0e;
      10'b1011001111: data <= 30'h391f4510;
      10'b1011010000: data <= 30'h392a9642;
      10'b1011010001: data <= 30'h3935dea4;
      10'b1011010010: data <= 30'h39411e33;
      10'b1011010011: data <= 30'h394c54ee;
      10'b1011010100: data <= 30'h395782d3;
      10'b1011010101: data <= 30'h3962a7e0;
      10'b1011010110: data <= 30'h396dc414;
      10'b1011010111: data <= 30'h3978d76c;
      10'b1011011000: data <= 30'h3983e1e8;
      10'b1011011001: data <= 30'h398ee385;
      10'b1011011010: data <= 30'h3999dc42;
      10'b1011011011: data <= 30'h39a4cc1c;
      10'b1011011100: data <= 30'h39afb313;
      10'b1011011101: data <= 30'h39ba9125;
      10'b1011011110: data <= 30'h39c5664f;
      10'b1011011111: data <= 30'h39d03291;
      10'b1011100000: data <= 30'h39daf5e8;
      10'b1011100001: data <= 30'h39e5b054;
      10'b1011100010: data <= 30'h39f061d2;
      10'b1011100011: data <= 30'h39fb0a60;
      10'b1011100100: data <= 30'h3a05a9fd;
      10'b1011100101: data <= 30'h3a1040a8;
      10'b1011100110: data <= 30'h3a1ace5f;
      10'b1011100111: data <= 30'h3a25531f;
      10'b1011101000: data <= 30'h3a2fcee8;
      10'b1011101001: data <= 30'h3a3a41b9;
      10'b1011101010: data <= 30'h3a44ab8e;
      10'b1011101011: data <= 30'h3a4f0c67;
      10'b1011101100: data <= 30'h3a596442;
      10'b1011101101: data <= 30'h3a63b31d;
      10'b1011101110: data <= 30'h3a6df8f8;
      10'b1011101111: data <= 30'h3a7835cf;
      10'b1011110000: data <= 30'h3a8269a3;
      10'b1011110001: data <= 30'h3a8c9470;
      10'b1011110010: data <= 30'h3a96b636;
      10'b1011110011: data <= 30'h3aa0cef3;
      10'b1011110100: data <= 30'h3aaadea6;
      10'b1011110101: data <= 30'h3ab4e54c;
      10'b1011110110: data <= 30'h3abee2e5;
      10'b1011110111: data <= 30'h3ac8d76f;
      10'b1011111000: data <= 30'h3ad2c2e8;
      10'b1011111001: data <= 30'h3adca54e;
      10'b1011111010: data <= 30'h3ae67ea1;
      10'b1011111011: data <= 30'h3af04edf;
      10'b1011111100: data <= 30'h3afa1605;
      10'b1011111101: data <= 30'h3b03d414;
      10'b1011111110: data <= 30'h3b0d8909;
      10'b1011111111: data <= 30'h3b1734e2;
      10'b1100000000: data <= 30'h3b20d79e;
      10'b1100000001: data <= 30'h3b2a713d;
      10'b1100000010: data <= 30'h3b3401bb;
      10'b1100000011: data <= 30'h3b3d8918;
      10'b1100000100: data <= 30'h3b470753;
      10'b1100000101: data <= 30'h3b507c69;
      10'b1100000110: data <= 30'h3b59e85a;
      10'b1100000111: data <= 30'h3b634b23;
      10'b1100001000: data <= 30'h3b6ca4c4;
      10'b1100001001: data <= 30'h3b75f53c;
      10'b1100001010: data <= 30'h3b7f3c87;
      10'b1100001011: data <= 30'h3b887aa6;
      10'b1100001100: data <= 30'h3b91af97;
      10'b1100001101: data <= 30'h3b9adb57;
      10'b1100001110: data <= 30'h3ba3fde7;
      10'b1100001111: data <= 30'h3bad1744;
      10'b1100010000: data <= 30'h3bb6276e;
      10'b1100010001: data <= 30'h3bbf2e62;
      10'b1100010010: data <= 30'h3bc82c1f;
      10'b1100010011: data <= 30'h3bd120a4;
      10'b1100010100: data <= 30'h3bda0bf0;
      10'b1100010101: data <= 30'h3be2ee01;
      10'b1100010110: data <= 30'h3bebc6d5;
      10'b1100010111: data <= 30'h3bf4966c;
      10'b1100011000: data <= 30'h3bfd5cc4;
      10'b1100011001: data <= 30'h3c0619dc;
      10'b1100011010: data <= 30'h3c0ecdb2;
      10'b1100011011: data <= 30'h3c177845;
      10'b1100011100: data <= 30'h3c201994;
      10'b1100011101: data <= 30'h3c28b19e;
      10'b1100011110: data <= 30'h3c314060;
      10'b1100011111: data <= 30'h3c39c5da;
      10'b1100100000: data <= 30'h3c42420a;
      10'b1100100001: data <= 30'h3c4ab4ef;
      10'b1100100010: data <= 30'h3c531e88;
      10'b1100100011: data <= 30'h3c5b7ed4;
      10'b1100100100: data <= 30'h3c63d5d1;
      10'b1100100101: data <= 30'h3c6c237e;
      10'b1100100110: data <= 30'h3c7467d9;
      10'b1100100111: data <= 30'h3c7ca2e2;
      10'b1100101000: data <= 30'h3c84d496;
      10'b1100101001: data <= 30'h3c8cfcf6;
      10'b1100101010: data <= 30'h3c951bff;
      10'b1100101011: data <= 30'h3c9d31b0;
      10'b1100101100: data <= 30'h3ca53e09;
      10'b1100101101: data <= 30'h3cad4107;
      10'b1100101110: data <= 30'h3cb53aaa;
      10'b1100101111: data <= 30'h3cbd2af0;
      10'b1100110000: data <= 30'h3cc511d9;
      10'b1100110001: data <= 30'h3cccef62;
      10'b1100110010: data <= 30'h3cd4c38b;
      10'b1100110011: data <= 30'h3cdc8e52;
      10'b1100110100: data <= 30'h3ce44fb7;
      10'b1100110101: data <= 30'h3cec07b8;
      10'b1100110110: data <= 30'h3cf3b653;
      10'b1100110111: data <= 30'h3cfb5b89;
      10'b1100111000: data <= 30'h3d02f757;
      10'b1100111001: data <= 30'h3d0a89bc;
      10'b1100111010: data <= 30'h3d1212b7;
      10'b1100111011: data <= 30'h3d199248;
      10'b1100111100: data <= 30'h3d21086c;
      10'b1100111101: data <= 30'h3d287523;
      10'b1100111110: data <= 30'h3d2fd86c;
      10'b1100111111: data <= 30'h3d373245;
      10'b1101000000: data <= 30'h3d3e82ae;
      10'b1101000001: data <= 30'h3d45c9a4;
      10'b1101000010: data <= 30'h3d4d0728;
      10'b1101000011: data <= 30'h3d543b37;
      10'b1101000100: data <= 30'h3d5b65d2;
      10'b1101000101: data <= 30'h3d6286f6;
      10'b1101000110: data <= 30'h3d699ea3;
      10'b1101000111: data <= 30'h3d70acd7;
      10'b1101001000: data <= 30'h3d77b192;
      10'b1101001001: data <= 30'h3d7eacd2;
      10'b1101001010: data <= 30'h3d859e96;
      10'b1101001011: data <= 30'h3d8c86de;
      10'b1101001100: data <= 30'h3d9365a8;
      10'b1101001101: data <= 30'h3d9a3af2;
      10'b1101001110: data <= 30'h3da106bd;
      10'b1101001111: data <= 30'h3da7c907;
      10'b1101010000: data <= 30'h3dae81cf;
      10'b1101010001: data <= 30'h3db53113;
      10'b1101010010: data <= 30'h3dbbd6d4;
      10'b1101010011: data <= 30'h3dc2730f;
      10'b1101010100: data <= 30'h3dc905c5;
      10'b1101010101: data <= 30'h3dcf8ef3;
      10'b1101010110: data <= 30'h3dd60e99;
      10'b1101010111: data <= 30'h3ddc84b5;
      10'b1101011000: data <= 30'h3de2f148;
      10'b1101011001: data <= 30'h3de9544f;
      10'b1101011010: data <= 30'h3defadca;
      10'b1101011011: data <= 30'h3df5fdb8;
      10'b1101011100: data <= 30'h3dfc4418;
      10'b1101011101: data <= 30'h3e0280e9;
      10'b1101011110: data <= 30'h3e08b42a;
      10'b1101011111: data <= 30'h3e0eddd9;
      10'b1101100000: data <= 30'h3e14fdf7;
      10'b1101100001: data <= 30'h3e1b1482;
      10'b1101100010: data <= 30'h3e212179;
      10'b1101100011: data <= 30'h3e2724db;
      10'b1101100100: data <= 30'h3e2d1ea8;
      10'b1101100101: data <= 30'h3e330ede;
      10'b1101100110: data <= 30'h3e38f57c;
      10'b1101100111: data <= 30'h3e3ed282;
      10'b1101101000: data <= 30'h3e44a5ef;
      10'b1101101001: data <= 30'h3e4a6fc1;
      10'b1101101010: data <= 30'h3e502ff9;
      10'b1101101011: data <= 30'h3e55e694;
      10'b1101101100: data <= 30'h3e5b9392;
      10'b1101101101: data <= 30'h3e6136f3;
      10'b1101101110: data <= 30'h3e66d0b4;
      10'b1101101111: data <= 30'h3e6c60d7;
      10'b1101110000: data <= 30'h3e71e759;
      10'b1101110001: data <= 30'h3e77643a;
      10'b1101110010: data <= 30'h3e7cd778;
      10'b1101110011: data <= 30'h3e824114;
      10'b1101110100: data <= 30'h3e87a10c;
      10'b1101110101: data <= 30'h3e8cf75f;
      10'b1101110110: data <= 30'h3e92440d;
      10'b1101110111: data <= 30'h3e978715;
      10'b1101111000: data <= 30'h3e9cc076;
      10'b1101111001: data <= 30'h3ea1f02f;
      10'b1101111010: data <= 30'h3ea7163f;
      10'b1101111011: data <= 30'h3eac32a6;
      10'b1101111100: data <= 30'h3eb14563;
      10'b1101111101: data <= 30'h3eb64e75;
      10'b1101111110: data <= 30'h3ebb4ddb;
      10'b1101111111: data <= 30'h3ec04394;
      10'b1110000000: data <= 30'h3ec52fa0;
      10'b1110000001: data <= 30'h3eca11fe;
      10'b1110000010: data <= 30'h3eceeaad;
      10'b1110000011: data <= 30'h3ed3b9ad;
      10'b1110000100: data <= 30'h3ed87efc;
      10'b1110000101: data <= 30'h3edd3a9a;
      10'b1110000110: data <= 30'h3ee1ec87;
      10'b1110000111: data <= 30'h3ee694c1;
      10'b1110001000: data <= 30'h3eeb3347;
      10'b1110001001: data <= 30'h3eefc81a;
      10'b1110001010: data <= 30'h3ef45338;
      10'b1110001011: data <= 30'h3ef8d4a1;
      10'b1110001100: data <= 30'h3efd4c54;
      10'b1110001101: data <= 30'h3f01ba50;
      10'b1110001110: data <= 30'h3f061e95;
      10'b1110001111: data <= 30'h3f0a7921;
      10'b1110010000: data <= 30'h3f0ec9f5;
      10'b1110010001: data <= 30'h3f13110f;
      10'b1110010010: data <= 30'h3f174e70;
      10'b1110010011: data <= 30'h3f1b8215;
      10'b1110010100: data <= 30'h3f1fabff;
      10'b1110010101: data <= 30'h3f23cc2e;
      10'b1110010110: data <= 30'h3f27e29f;
      10'b1110010111: data <= 30'h3f2bef53;
      10'b1110011000: data <= 30'h3f2ff24a;
      10'b1110011001: data <= 30'h3f33eb81;
      10'b1110011010: data <= 30'h3f37dafa;
      10'b1110011011: data <= 30'h3f3bc0b3;
      10'b1110011100: data <= 30'h3f3f9cab;
      10'b1110011101: data <= 30'h3f436ee3;
      10'b1110011110: data <= 30'h3f473759;
      10'b1110011111: data <= 30'h3f4af60d;
      10'b1110100000: data <= 30'h3f4eaafe;
      10'b1110100001: data <= 30'h3f52562c;
      10'b1110100010: data <= 30'h3f55f796;
      10'b1110100011: data <= 30'h3f598f3c;
      10'b1110100100: data <= 30'h3f5d1d1d;
      10'b1110100101: data <= 30'h3f60a138;
      10'b1110100110: data <= 30'h3f641b8d;
      10'b1110100111: data <= 30'h3f678c1c;
      10'b1110101000: data <= 30'h3f6af2e3;
      10'b1110101001: data <= 30'h3f6e4fe3;
      10'b1110101010: data <= 30'h3f71a31b;
      10'b1110101011: data <= 30'h3f74ec8a;
      10'b1110101100: data <= 30'h3f782c30;
      10'b1110101101: data <= 30'h3f7b620c;
      10'b1110101110: data <= 30'h3f7e8e1e;
      10'b1110101111: data <= 30'h3f81b065;
      10'b1110110000: data <= 30'h3f84c8e2;
      10'b1110110001: data <= 30'h3f87d792;
      10'b1110110010: data <= 30'h3f8adc77;
      10'b1110110011: data <= 30'h3f8dd78f;
      10'b1110110100: data <= 30'h3f90c8da;
      10'b1110110101: data <= 30'h3f93b058;
      10'b1110110110: data <= 30'h3f968e07;
      10'b1110110111: data <= 30'h3f9961e8;
      10'b1110111000: data <= 30'h3f9c2bfb;
      10'b1110111001: data <= 30'h3f9eec3e;
      10'b1110111010: data <= 30'h3fa1a2b2;
      10'b1110111011: data <= 30'h3fa44f55;
      10'b1110111100: data <= 30'h3fa6f228;
      10'b1110111101: data <= 30'h3fa98b2a;
      10'b1110111110: data <= 30'h3fac1a5b;
      10'b1110111111: data <= 30'h3fae9fbb;
      10'b1111000000: data <= 30'h3fb11b48;
      10'b1111000001: data <= 30'h3fb38d02;
      10'b1111000010: data <= 30'h3fb5f4ea;
      10'b1111000011: data <= 30'h3fb852ff;
      10'b1111000100: data <= 30'h3fbaa740;
      10'b1111000101: data <= 30'h3fbcf1ad;
      10'b1111000110: data <= 30'h3fbf3246;
      10'b1111000111: data <= 30'h3fc1690a;
      10'b1111001000: data <= 30'h3fc395f9;
      10'b1111001001: data <= 30'h3fc5b913;
      10'b1111001010: data <= 30'h3fc7d258;
      10'b1111001011: data <= 30'h3fc9e1c6;
      10'b1111001100: data <= 30'h3fcbe75e;
      10'b1111001101: data <= 30'h3fcde320;
      10'b1111001110: data <= 30'h3fcfd50b;
      10'b1111001111: data <= 30'h3fd1bd1e;
      10'b1111010000: data <= 30'h3fd39b5a;
      10'b1111010001: data <= 30'h3fd56fbe;
      10'b1111010010: data <= 30'h3fd73a4a;
      10'b1111010011: data <= 30'h3fd8fafe;
      10'b1111010100: data <= 30'h3fdab1d9;
      10'b1111010101: data <= 30'h3fdc5edc;
      10'b1111010110: data <= 30'h3fde0205;
      10'b1111010111: data <= 30'h3fdf9b55;
      10'b1111011000: data <= 30'h3fe12acb;
      10'b1111011001: data <= 30'h3fe2b067;
      10'b1111011010: data <= 30'h3fe42c2a;
      10'b1111011011: data <= 30'h3fe59e12;
      10'b1111011100: data <= 30'h3fe7061f;
      10'b1111011101: data <= 30'h3fe86452;
      10'b1111011110: data <= 30'h3fe9b8a9;
      10'b1111011111: data <= 30'h3feb0326;
      10'b1111100000: data <= 30'h3fec43c7;
      10'b1111100001: data <= 30'h3fed7a8c;
      10'b1111100010: data <= 30'h3feea776;
      10'b1111100011: data <= 30'h3fefca84;
      10'b1111100100: data <= 30'h3ff0e3b6;
      10'b1111100101: data <= 30'h3ff1f30b;
      10'b1111100110: data <= 30'h3ff2f884;
      10'b1111100111: data <= 30'h3ff3f420;
      10'b1111101000: data <= 30'h3ff4e5e0;
      10'b1111101001: data <= 30'h3ff5cdc3;
      10'b1111101010: data <= 30'h3ff6abc8;
      10'b1111101011: data <= 30'h3ff77ff1;
      10'b1111101100: data <= 30'h3ff84a3c;
      10'b1111101101: data <= 30'h3ff90aaa;
      10'b1111101110: data <= 30'h3ff9c13a;
      10'b1111101111: data <= 30'h3ffa6dec;
      10'b1111110000: data <= 30'h3ffb10c1;
      10'b1111110001: data <= 30'h3ffba9b8;
      10'b1111110010: data <= 30'h3ffc38d1;
      10'b1111110011: data <= 30'h3ffcbe0c;
      10'b1111110100: data <= 30'h3ffd3969;
      10'b1111110101: data <= 30'h3ffdaae7;
      10'b1111110110: data <= 30'h3ffe1288;
      10'b1111110111: data <= 30'h3ffe704a;
      10'b1111111000: data <= 30'h3ffec42d;
      10'b1111111001: data <= 30'h3fff0e32;
      10'b1111111010: data <= 30'h3fff4e59;
      10'b1111111011: data <= 30'h3fff84a1;
      10'b1111111100: data <= 30'h3fffb10b;
      10'b1111111101: data <= 30'h3fffd396;
      10'b1111111110: data <= 30'h3fffec43;
      10'b1111111111: data <= 30'h3ffffb11;

      default: data <= 30'h0;
    endcase
  end
endmodule
     